module generator;
endmodule // generator
