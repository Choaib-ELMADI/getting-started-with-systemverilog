class generator;
endclass // generator
