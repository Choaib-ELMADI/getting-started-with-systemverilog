class driver extends uvm_driver;
    function new();
    endfunction // new

endclass // driver
