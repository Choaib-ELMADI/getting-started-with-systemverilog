class class_name;
    bit [7:0] bus;
    int       range;

    function function_name;
    endfunction // function_name

    task task_name;
    endtask // task_name

endclass // class_name
