module test;
endmodule // test
