class monitor extends uvm_monitor;
    function new();
    endfunction // new

endclass // monitor
