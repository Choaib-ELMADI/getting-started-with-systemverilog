interface full_adder_if;

    // Signals
    logic a, b, c_in;
    logic s, c_out;

    // Clocking block

    // Modport

endinterface // full_adder_if
