class scoreboard extends uvm_scoreboard;
    bit [7:0] mem [0:3];

    function new();
    endfunction // new

endclass // scoreboard
