`include "generator.sv"
`include "full_adder_if.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"

class environment;
    generator  gen;
    driver     drv;
    monitor    mnt;
    scoreboard scb;

    mailbox gen2drv;
    mailbox mnt2scb;

    virtual full_adder_if vir_interface_inst;

    function new(virtual full_adder_if vir_interface_inst);
        this.vir_interface_inst = vir_interface_inst;

        gen2drv = new();
        mnt2scb = new();

        gen = new(gen2drv);
        drv = new();
        mnt = new();
        scb = new();

        drv.vir_interface_inst = vir_interface_inst;
        drv.gen2drv = gen2drv;

        mnt.vir_interface_inst = vir_interface_inst;
        mnt.mnt2scb = mnt2scb;

        scb.mnt2scb = mnt2scb;
    endfunction // new

    task test_run();
        fork
            gen.main();
            drv.main();
            mnt.main();
            scb.main();
        join
    endtask // test_run

endclass // environment
