interface interface_;

    // Signals
    logic a, b, c_in;
    logic s, c_out;

    // Clocking block

    // Modport

endinterface // interface_
