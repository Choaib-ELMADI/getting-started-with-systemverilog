class scoreboard;
    mailbox mnt2scb;

    // Local memory
    bit [7:0] mem [0:3];

    function new();
    endfunction // new

endclass // scoreboard
