module interface_;
endmodule // interface_
