class monitor;
    mailbox mnt2scb;

    function new();
    endfunction // new

endclass // monitor
