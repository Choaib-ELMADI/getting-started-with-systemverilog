class driver;
    mailbox gen2drv;

    function new();
    endfunction // new

endclass // driver
